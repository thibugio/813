library verilog;
use verilog.vl_types.all;
entity testfifo is
end testfifo;
