/* testssp.v
    testbench for ssp module
*/

module testssp;

endmodule
