library verilog;
use verilog.vl_types.all;
entity testStructural is
end testStructural;
